GLOBAL
gameDifficulty:MEDIUM
SUSPECTS
classSuspect:Innocent
fullNameSuspect:Antoine Fourmond
ageSuspect     :42
sexSuspect     :homme
lookSuspect    :look1
aspectSuspect  :aspect2
stressSuspect     :69
cooperationSuspect:51
innocentSuspect   :false
alibiSuspect:alibi-false
seenSuspect :J'ai vu vu-false
heardSuspect:j'ai entendu entendu-false
classSuspect:Murderer
fullNameSuspect:Claire Juzeau
ageSuspect     :79
sexSuspect     :femme
lookSuspect    :look2
aspectSuspect  :aspect2
stressSuspect     :61
cooperationSuspect:0
innocentSuspect   :false
alibiSuspect:null
seenSuspect :null
heardSuspect:null
motiveMurderer:la folie
classSuspect:Innocent
fullNameSuspect:Pierre Boore
ageSuspect     :52
sexSuspect     :homme
lookSuspect    :look1
aspectSuspect  :aspect2
stressSuspect     :58
cooperationSuspect:67
innocentSuspect   :false
alibiSuspect:alibi-false
seenSuspect :J'ai vu vu-false
heardSuspect:j'ai entendu entendu-false
classSuspect:Innocent
fullNameSuspect:Jean Deolivera
ageSuspect     :57
sexSuspect     :homme
lookSuspect    :look2
aspectSuspect  :aspect2
stressSuspect     :58
cooperationSuspect:44
innocentSuspect   :false
alibiSuspect:alibi-false
seenSuspect :J'ai vu vu-false
heardSuspect:j'ai entendu entendu-false
classSuspect:CrimePartner
fullNameSuspect:Luc Pasquier
ageSuspect     :69
sexSuspect     :homme
lookSuspect    :look1
aspectSuspect  :aspect1
stressSuspect     :40
cooperationSuspect:49
innocentSuspect   :false
alibiSuspect:alibi-false
seenSuspect :null
heardSuspect:null
classSuspect:Innocent
fullNameSuspect:Laure Deolivera
ageSuspect     :52
sexSuspect     :femme
lookSuspect    :look1
aspectSuspect  :aspect2
stressSuspect     :40
cooperationSuspect:40
innocentSuspect   :false
alibiSuspect:alibi-false
seenSuspect :J'ai vu vu-false
heardSuspect:j'ai entendu entendu-false
classSuspect:Innocent
fullNameSuspect:Alexandre Deolivera
ageSuspect     :36
sexSuspect     :homme
lookSuspect    :look1
aspectSuspect  :aspect2
stressSuspect     :51
cooperationSuspect:45
innocentSuspect   :false
alibiSuspect:alibi-false
seenSuspect :J'ai vu vu-false
heardSuspect:j'ai entendu entendu-false
classSuspect:Innocent
fullNameSuspect:Antoine Juzeau
ageSuspect     :20
sexSuspect     :homme
lookSuspect    :look2
aspectSuspect  :aspect1
stressSuspect     :46
cooperationSuspect:55
innocentSuspect   :false
alibiSuspect:alibi-false
seenSuspect :J'ai vu vu-false
heardSuspect:j'ai entendu entendu-false
classSuspect:Innocent
fullNameSuspect:Jean Bomy
ageSuspect     :29
sexSuspect     :homme
lookSuspect    :look1
aspectSuspect  :aspect2
stressSuspect     :48
cooperationSuspect:66
innocentSuspect   :false
alibiSuspect:alibi-false
seenSuspect :J'ai vu vu-false
heardSuspect:j'ai entendu entendu-false
classSuspect:Innocent
fullNameSuspect:Alexandre Bomy
ageSuspect     :31
sexSuspect     :homme
lookSuspect    :look1
aspectSuspect  :aspect2
stressSuspect     :57
cooperationSuspect:45
innocentSuspect   :false
alibiSuspect:alibi-false
seenSuspect :J'ai vu vu-false
heardSuspect:j'ai entendu entendu-false
classSuspect:Innocent
fullNameSuspect:Jean Pasquier
ageSuspect     :60
sexSuspect     :homme
lookSuspect    :look2
aspectSuspect  :aspect1
stressSuspect     :67
cooperationSuspect:40
innocentSuspect   :false
alibiSuspect:alibi-false
seenSuspect :J'ai vu vu-false
heardSuspect:j'ai entendu entendu-false
classSuspect:Innocent
fullNameSuspect:Paul Boore
ageSuspect     :59
sexSuspect     :homme
lookSuspect    :look1
aspectSuspect  :aspect2
stressSuspect     :56
cooperationSuspect:40
innocentSuspect   :false
alibiSuspect:alibi-false
seenSuspect :J'ai vu vu-false
heardSuspect:j'ai entendu entendu-false
VICTIM
fullNameVictim:Antoine Juzeau
sexVictim     :homme
ageVictim     :53
deathDateVictim :il y a 6 jours, à 19h15
deathCauseVictim:blessure par balle
VICTIMPROOF
contentProofVictim:contenu
WEAPON
typeWeapon:type d'arme
WEAPONPROOF
contentProofWeapon:contenu
contentProofWeapon:contenu
SCENE
typeScene:type d'endroit
SCENEPROOF
contentProofScene:contenu
contentProofScene:contenu
INVESTIGATOR
nameInvestigator:Thib Juzeau
SexInvestigator:homme
manipulationInvestigator:52
intelligenceInvestigator:52
supposedMurderer:null
supposedVictim  :null
supposedWeapon  :null
supposedMobile  :null
CLUES
