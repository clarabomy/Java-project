fileName : fullName
gameDifficulty : SIMPLE
SexInvestigator : homme
manipulationInvestigator : 60
intelligenceInvestigator : 75
supposedMurderer : null
supposedVictim   : null
supposedWeapon   : null
supposedMobile   : null
classSuspect : Innocent
fullNameSuspect : prenom innocent1
ageSuspect      : 35
sexSuspect      : homme
lookSuspect     : look
aspectSuspect   : aspect physique
stressSuspect      : 50
cooperationSuspect : 30
innocentSuspect    : false
alibiContentSuspect : alibi
alibiSuspectIsLie   : false
seenContentSuspect  : J'ai vu vu
seenSuspectIsLie    : false
heardContentSuspect : j'ai entendu entendu
heardSuspectIsLie   : false
classSuspect : Innocent
fullNameSuspect : prenom innocent3
ageSuspect      : 35
sexSuspect      : homme
lookSuspect     : look
aspectSuspect   : aspect physique
stressSuspect      : 50
cooperationSuspect : 30
innocentSuspect    : false
alibiContentSuspect : alibi
alibiSuspectIsLie   : false
seenContentSuspect  : J'ai vu vu
seenSuspectIsLie    : false
heardContentSuspect : j'ai entendu entendu
heardSuspectIsLie   : false
classSuspect : Murderer
fullNameSuspect : prenom criminel
ageSuspect      : 35
sexSuspect      : homme
lookSuspect     : look
aspectSuspect   : aspect physique
stressSuspect      : 50
cooperationSuspect : 0
innocentSuspect    : false
alibiContentSuspect : null
alibiSuspectIsLie   : null
seenContentSuspect  : null
seenSuspectIsLie    : null
heardContentSuspect : null
heardSuspectIsLie   : null
motiveMurderer : motivation
classSuspect : CrimePartner
fullNameSuspect : prenom partner
ageSuspect      : 35
sexSuspect      : homme
lookSuspect     : look
aspectSuspect   : aspect physique
stressSuspect      : 50
cooperationSuspect : 30
innocentSuspect    : false
alibiContentSuspect : alibi
alibiSuspectIsLie   : false
seenContentSuspect  : null
seenSuspectIsLie    : null
heardContentSuspect : null
heardSuspectIsLie   : null
classSuspect : Innocent
fullNameSuspect : prenom innocent2
ageSuspect      : 35
sexSuspect      : homme
lookSuspect     : look
aspectSuspect   : aspect physique
stressSuspect      : 50
cooperationSuspect : 30
innocentSuspect    : false
alibiContentSuspect : alibi
alibiSuspectIsLie   : false
seenContentSuspect  : J'ai vu vu
seenSuspectIsLie    : false
heardContentSuspect : j'ai entendu entendu
heardSuspectIsLie   : false
classSuspect : Innocent
fullNameSuspect : prenom innocent0
ageSuspect      : 35
sexSuspect      : homme
lookSuspect     : look
aspectSuspect   : aspect physique
stressSuspect      : 50
cooperationSuspect : 30
innocentSuspect    : false
alibiContentSuspect : alibi
alibiSuspectIsLie   : false
seenContentSuspect  : J'ai vu vu
seenSuspectIsLie    : false
heardContentSuspect : j'ai entendu entendu
heardSuspectIsLie   : false
fullNameVictim : Prenom Nom
sexVictim      : homme
ageVictim      : 35
deathDateVictim  : date et heure de la mort
deathCauseVictim : cause de la mort
contentProofVictim : contenu
typeWeapon : type d'arme
contentProofWeapon : contenu
typeScene : type d'endroit
contentProofScene : contenu
